module comparator4bit(a,b,eq,gr,le);
input [3:0]a,b;
output reg eq,gr,le;
always @(a,b)
begin
if (a==b)
begin
eq=1;le=0;gr=0;
end
else if (a<b)
begin
eq=0;le=1;gr=0;
end
else
begin
eq=0;le=0;gr=1;
end
end
endmodule
