module Ad_sub_4bit(a,b,sel,CB,r);  ///when sel=1 thn it performs subtraction else addition///
input [3:0]a;
input [3:0]b;
input sel;
output [3:0]r;
output CB;
wire [3:0]w;
wire [2:0]cr;

xor f1(b[0],sel,w[0]);
full_adder fa1(w[0],a[0],sel,cr[0],r[0]);

xor f2(b[1],sel,w[1]);
full_adder fa2(w[1],a[1],cr[0],cr[1],r[1]);

xor f3(b[2],sel,w[2]);
full_adder fa3(w[2],a[2],cr[1],cr[2],r[2]);

xor f4(b[3],sel,w[3]);
full_adder fa4(w[3],a[3],cr[2],CB,r[3]);

endmodule
 

////full adder/////
module full_adder(X,Y,Z,C,S);
input X,Y,Z;
output C,S;
assign S=X^Y^Z;
assign C=(X&(Y^Z))|(Y&Z);
endmodule
