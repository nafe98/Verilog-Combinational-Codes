module ALU(A,B,S,Y);
input [1:0]A,B,S;
output reg [1:0]Y;

always@*
begin
case(S)
2'b00:Y=A+B;
2'b01:Y=A&B;
2'b10:Y=A|B;
2'b11:Y=A^B;
endcase
end
endmodule
